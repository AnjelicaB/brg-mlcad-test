//========================================================================
// Prob06p06_comb_codes_penc_16to4_ref
//========================================================================
// SPDX-License-Identifier: MIT
// Author : Christopher Batten, NVIDIA
// Date   : May 20, 2024

module RefModule
(
  input  logic [15:0] in_,
  output logic [ 3:0] out
);

  always @(*) begin
    casez ( in_ )

      16'b????_????_????_???1 : out = 4'd0;
      16'b????_????_????_??10 : out = 4'd1;
      16'b????_????_????_?100 : out = 4'd2;
      16'b????_????_????_1000 : out = 4'd3;

      16'b????_????_???1_0000 : out = 4'd4;
      16'b????_????_??10_0000 : out = 4'd5;
      16'b????_????_?100_0000 : out = 4'd6;
      16'b????_????_1000_0000 : out = 4'd7;

      16'b????_???1_0000_0000 : out = 4'd8;
      16'b????_??10_0000_0000 : out = 4'd9;
      16'b????_?100_0000_0000 : out = 4'd10;
      16'b????_1000_0000_0000 : out = 4'd11;

      16'b???1_0000_0000_0000 : out = 4'd12;
      16'b??10_0000_0000_0000 : out = 4'd13;
      16'b?100_0000_0000_0000 : out = 4'd14;
      16'b1000_0000_0000_0000 : out = 4'd15;

      default                 : out = 4'd0;

    endcase
  end

endmodule

