//========================================================================
// Prob01p04_comb_const_32b_value_ref
//========================================================================
// SPDX-License-Identifier: MIT
// Author : Christopher Batten, NVIDIA
// Date   : May 20, 2024

module RefModule
(
  output logic [31:0] out
);

  assign out = 32'hdeadbeef;

endmodule

