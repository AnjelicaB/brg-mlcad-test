//========================================================================
// Prob01p01_comb_const_zero_ref
//========================================================================
// SPDX-License-Identifier: MIT
// Author : Christopher Batten, NVIDIA
// Date   : May 20, 2024

module RefModule
(
  output logic zero
);

  assign zero = 1'b0;

endmodule

