//========================================================================
// Prob01p02_comb_const_one_ref
//========================================================================
// SPDX-License-Identifier: MIT
// Author : Christopher Batten, NVIDIA
// Date   : May 20, 2024

module RefModule
(
  output logic out
);

  assign out = 1'b1;

endmodule

