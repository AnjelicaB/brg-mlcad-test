//========================================================================
// Prob06p04_comb_codes_dec_4to16_ref
//========================================================================
// SPDX-License-Identifier: MIT
// Author : Christopher Batten, NVIDIA
// Date   : May 20, 2024

module RefModule
(
  input  logic [ 3:0] in_,
  output logic [15:0] out
);

  always @(*) begin
    case ( in_ )

      4'd0  : out = 16'b0000_0000_0000_0001;
      4'd1  : out = 16'b0000_0000_0000_0010;
      4'd2  : out = 16'b0000_0000_0000_0100;
      4'd3  : out = 16'b0000_0000_0000_1000;

      4'd4  : out = 16'b0000_0000_0001_0000;
      4'd5  : out = 16'b0000_0000_0010_0000;
      4'd6  : out = 16'b0000_0000_0100_0000;
      4'd7  : out = 16'b0000_0000_1000_0000;

      4'd8  : out = 16'b0000_0001_0000_0000;
      4'd9  : out = 16'b0000_0010_0000_0000;
      4'd10 : out = 16'b0000_0100_0000_0000;
      4'd11 : out = 16'b0000_1000_0000_0000;

      4'd12 : out = 16'b0001_0000_0000_0000;
      4'd13 : out = 16'b0010_0000_0000_0000;
      4'd14 : out = 16'b0100_0000_0000_0000;
      4'd15 : out = 16'b1000_0000_0000_0000;

    endcase
  end

endmodule

