//========================================================================
// Prob01p03_comb_const_lohi_ref
//========================================================================
// SPDX-License-Identifier: MIT
// Author : Christopher Batten, NVIDIA
// Date   : May 20, 2024

module RefModule
(
  output logic lo,
  output logic hi
);

  assign lo = 1'b0;
  assign hi = 1'b1;

endmodule

